`timescale 1 ps/ 1 psmodule blokus_fifo_tb;reg reset, clk, wr;reg [7:0] data_in;wire [7:0] data_out;blokus_fifo blokus_fifo_unit(.reset(reset), .clk(clk), .wr(wr), .data_in(data_in), .data_out(data_out));initial$monitor($time, " input = %h, output = %h", data_in, data_out);initialbegin reset = 0; clk = 0; wr = 0; data_in = 0; #3 reset = 1; #2 reset = 0;  #10 data_in = 8'h30; #2 wr = 1; #2 wr = 0; #10 data_in = 8'h32; #2 wr = 1; #2 wr = 0; #10 data_in = 8'h35; #2 wr = 1; #2 wr = 0; #1000 data_in = 8'h33; #2 wr = 1; #2 wr = 0; #100 data_in = 8'h61; #2 wr = 1; #2 wr = 0; #100 data_in = 8'h38; #2 wr = 1; #2 wr = 0; #100 data_in = 8'h71; #2 wr = 1; #2 wr = 0; #100 data_in = 8'h32; #2 wr = 1; #2 wr = 0;endalways	#1 clk = ~clk;initial	#1000 $finish;endmodule