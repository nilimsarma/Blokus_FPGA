`timescale 1 ns / 1 psmodule blokus_fifo_tb;reg reset, clk, wr, rd;reg [7:0] data_in;wire [7:0] data_out;blokus_fifo blokus_fifo_unit(.reset(reset), .clk(clk), .wr(wr), .rd(rd), .data_in(data_in), .data_out(data_out));initial $monitor($time, " input = %h, output = %h", data_in, data_out);initialbegin reset = 0; clk = 0; wr = 0; data_in = 0; #30 reset = 1; #40 reset = 0;  #100 data_in = 8'h30; #20 wr = 1; #20 wr = 0; #100 data_in = 8'h32; #20 wr = 1; #20 wr = 0; #100 data_in = 8'h35; #20 wr = 1; #20 wr = 0; #10000 data_in = 8'h33; #20 wr = 1; #20 wr = 0; #1000 data_in = 8'h61; #20 wr = 1; #20 wr = 0; #1000 data_in = 8'h38; #20 wr = 1; #20 wr = 0; #1000 data_in = 8'h71; #20 wr = 1; #20 wr = 0;  #1000 data_in = 8'h32; #20 wr = 1; #20 wr = 0;endalways	#10 clk = ~clk;initial	#10000 $finish;endmodule